module wave_rom(
	input clock,
	input [1:0] wave_select,
	input [7:0] phase,
	output [15:0] wave_out
	);

	wire [15:0] sine, saw, square;

	sine_rom s0 (clock, phase, sine);
	saw_rom s1 (clock, phase, saw);
	square_rom s2 (clock, phase, square);

	wave_mux u_wm(sine, saw, square, wave_select, wave_out);

endmodule

module wave_mux(
	input [15:0] sine, saw, square,
	input [1:0] wave_select,
	output reg [15:0] wave_out
	);

	always @ (*)
	begin
		case(wave_select)

		0: wave_out = sine;
		1: wave_out = saw;
		2: wave_out = square;

		default: wave_out = sine;

		endcase
	end

endmodule






//////////////////////////////////////////////////
////////////	Sin Wave ROM Table	//////////////
//////////////////////////////////////////////////
// produces a 2's comp, 16-bit, approximation
// of a sine wave, given an input phase (address)
module sine_rom (clock, address, sine);
input clock;
input [7:0] address;
output [15:0] sine;
reg signed [15:0] sine;
always@(posedge clock)
begin
    case(address)
    			8'h00: sine = 16'h0;
			8'h01: sine = 16'h324;
			8'h02: sine = 16'h647;
			8'h03: sine = 16'h96a;
			8'h04: sine = 16'hc8b;
			8'h05: sine = 16'hfab;
			8'h06: sine = 16'h12c7;
			8'h07: sine = 16'h15e1;
			8'h08: sine = 16'h18f8;
			8'h09: sine = 16'h1c0b;
			8'h0a: sine = 16'h1f19;
			8'h0b: sine = 16'h2223;
			8'h0c: sine = 16'h2527;
			8'h0d: sine = 16'h2826;
			8'h0e: sine = 16'h2b1e;
			8'h0f: sine = 16'h2e10;
			8'h10: sine = 16'h30fb;
			8'h11: sine = 16'h33de;
			8'h12: sine = 16'h36b9;
			8'h13: sine = 16'h398c;
			8'h14: sine = 16'h3c56;
			8'h15: sine = 16'h3f16;
			8'h16: sine = 16'h41cd;
			8'h17: sine = 16'h447a;
			8'h18: sine = 16'h471c;
			8'h19: sine = 16'h49b3;
			8'h1a: sine = 16'h4c3f;
			8'h1b: sine = 16'h4ebf;
			8'h1c: sine = 16'h5133;
			8'h1d: sine = 16'h539a;
			8'h1e: sine = 16'h55f4;
			8'h1f: sine = 16'h5842;
			8'h20: sine = 16'h5a81;
			8'h21: sine = 16'h5cb3;
			8'h22: sine = 16'h5ed6;
			8'h23: sine = 16'h60eb;
			8'h24: sine = 16'h62f1;
			8'h25: sine = 16'h64e7;
			8'h26: sine = 16'h66ce;
			8'h27: sine = 16'h68a5;
			8'h28: sine = 16'h6a6c;
			8'h29: sine = 16'h6c23;
			8'h2a: sine = 16'h6dc9;
			8'h2b: sine = 16'h6f5e;
			8'h2c: sine = 16'h70e1;
			8'h2d: sine = 16'h7254;
			8'h2e: sine = 16'h73b5;
			8'h2f: sine = 16'h7503;
			8'h30: sine = 16'h7640;
			8'h31: sine = 16'h776b;
			8'h32: sine = 16'h7883;
			8'h33: sine = 16'h7989;
			8'h34: sine = 16'h7a7c;
			8'h35: sine = 16'h7b5c;
			8'h36: sine = 16'h7c29;
			8'h37: sine = 16'h7ce2;
			8'h38: sine = 16'h7d89;
			8'h39: sine = 16'h7e1c;
			8'h3a: sine = 16'h7e9c;
			8'h3b: sine = 16'h7f08;
			8'h3c: sine = 16'h7f61;
			8'h3d: sine = 16'h7fa6;
			8'h3e: sine = 16'h7fd7;
			8'h3f: sine = 16'h7ff5;
			8'h40: sine = 16'h7fff;
			8'h41: sine = 16'h7ff5;
			8'h42: sine = 16'h7fd7;
			8'h43: sine = 16'h7fa6;
			8'h44: sine = 16'h7f61;
			8'h45: sine = 16'h7f08;
			8'h46: sine = 16'h7e9c;
			8'h47: sine = 16'h7e1c;
			8'h48: sine = 16'h7d89;
			8'h49: sine = 16'h7ce2;
			8'h4a: sine = 16'h7c29;
			8'h4b: sine = 16'h7b5c;
			8'h4c: sine = 16'h7a7c;
			8'h4d: sine = 16'h7989;
			8'h4e: sine = 16'h7883;
			8'h4f: sine = 16'h776b;
			8'h50: sine = 16'h7640;
			8'h51: sine = 16'h7503;
			8'h52: sine = 16'h73b5;
			8'h53: sine = 16'h7254;
			8'h54: sine = 16'h70e1;
			8'h55: sine = 16'h6f5e;
			8'h56: sine = 16'h6dc9;
			8'h57: sine = 16'h6c23;
			8'h58: sine = 16'h6a6c;
			8'h59: sine = 16'h68a5;
			8'h5a: sine = 16'h66ce;
			8'h5b: sine = 16'h64e7;
			8'h5c: sine = 16'h62f1;
			8'h5d: sine = 16'h60eb;
			8'h5e: sine = 16'h5ed6;
			8'h5f: sine = 16'h5cb3;
			8'h60: sine = 16'h5a81;
			8'h61: sine = 16'h5842;
			8'h62: sine = 16'h55f4;
			8'h63: sine = 16'h539a;
			8'h64: sine = 16'h5133;
			8'h65: sine = 16'h4ebf;
			8'h66: sine = 16'h4c3f;
			8'h67: sine = 16'h49b3;
			8'h68: sine = 16'h471c;
			8'h69: sine = 16'h447a;
			8'h6a: sine = 16'h41cd;
			8'h6b: sine = 16'h3f16;
			8'h6c: sine = 16'h3c56;
			8'h6d: sine = 16'h398c;
			8'h6e: sine = 16'h36b9;
			8'h6f: sine = 16'h33de;
			8'h70: sine = 16'h30fb;
			8'h71: sine = 16'h2e10;
			8'h72: sine = 16'h2b1e;
			8'h73: sine = 16'h2826;
			8'h74: sine = 16'h2527;
			8'h75: sine = 16'h2223;
			8'h76: sine = 16'h1f19;
			8'h77: sine = 16'h1c0b;
			8'h78: sine = 16'h18f8;
			8'h79: sine = 16'h15e1;
			8'h7a: sine = 16'h12c7;
			8'h7b: sine = 16'hfab;
			8'h7c: sine = 16'hc8b;
			8'h7d: sine = 16'h96a;
			8'h7e: sine = 16'h647;
			8'h7f: sine = 16'h324;
			8'h80: sine = 16'h0;
			8'h81: sine = 16'hfcdc;
			8'h82: sine = 16'hf9b9;
			8'h83: sine = 16'hf696;
			8'h84: sine = 16'hf375;
			8'h85: sine = 16'hf055;
			8'h86: sine = 16'hed39;
			8'h87: sine = 16'hea1f;
			8'h88: sine = 16'he708;
			8'h89: sine = 16'he3f5;
			8'h8a: sine = 16'he0e7;
			8'h8b: sine = 16'hdddd;
			8'h8c: sine = 16'hdad9;
			8'h8d: sine = 16'hd7da;
			8'h8e: sine = 16'hd4e2;
			8'h8f: sine = 16'hd1f0;
			8'h90: sine = 16'hcf05;
			8'h91: sine = 16'hcc22;
			8'h92: sine = 16'hc947;
			8'h93: sine = 16'hc674;
			8'h94: sine = 16'hc3aa;
			8'h95: sine = 16'hc0ea;
			8'h96: sine = 16'hbe33;
			8'h97: sine = 16'hbb86;
			8'h98: sine = 16'hb8e4;
			8'h99: sine = 16'hb64d;
			8'h9a: sine = 16'hb3c1;
			8'h9b: sine = 16'hb141;
			8'h9c: sine = 16'haecd;
			8'h9d: sine = 16'hac66;
			8'h9e: sine = 16'haa0c;
			8'h9f: sine = 16'ha7be;
			8'ha0: sine = 16'ha57f;
			8'ha1: sine = 16'ha34d;
			8'ha2: sine = 16'ha12a;
			8'ha3: sine = 16'h9f15;
			8'ha4: sine = 16'h9d0f;
			8'ha5: sine = 16'h9b19;
			8'ha6: sine = 16'h9932;
			8'ha7: sine = 16'h975b;
			8'ha8: sine = 16'h9594;
			8'ha9: sine = 16'h93dd;
			8'haa: sine = 16'h9237;
			8'hab: sine = 16'h90a2;
			8'hac: sine = 16'h8f1f;
			8'had: sine = 16'h8dac;
			8'hae: sine = 16'h8c4b;
			8'haf: sine = 16'h8afd;
			8'hb0: sine = 16'h89c0;
			8'hb1: sine = 16'h8895;
			8'hb2: sine = 16'h877d;
			8'hb3: sine = 16'h8677;
			8'hb4: sine = 16'h8584;
			8'hb5: sine = 16'h84a4;
			8'hb6: sine = 16'h83d7;
			8'hb7: sine = 16'h831e;
			8'hb8: sine = 16'h8277;
			8'hb9: sine = 16'h81e4;
			8'hba: sine = 16'h8164;
			8'hbb: sine = 16'h80f8;
			8'hbc: sine = 16'h809f;
			8'hbd: sine = 16'h805a;
			8'hbe: sine = 16'h8029;
			8'hbf: sine = 16'h800b;
			8'hc0: sine = 16'h8001;
			8'hc1: sine = 16'h800b;
			8'hc2: sine = 16'h8029;
			8'hc3: sine = 16'h805a;
			8'hc4: sine = 16'h809f;
			8'hc5: sine = 16'h80f8;
			8'hc6: sine = 16'h8164;
			8'hc7: sine = 16'h81e4;
			8'hc8: sine = 16'h8277;
			8'hc9: sine = 16'h831e;
			8'hca: sine = 16'h83d7;
			8'hcb: sine = 16'h84a4;
			8'hcc: sine = 16'h8584;
			8'hcd: sine = 16'h8677;
			8'hce: sine = 16'h877d;
			8'hcf: sine = 16'h8895;
			8'hd0: sine = 16'h89c0;
			8'hd1: sine = 16'h8afd;
			8'hd2: sine = 16'h8c4b;
			8'hd3: sine = 16'h8dac;
			8'hd4: sine = 16'h8f1f;
			8'hd5: sine = 16'h90a2;
			8'hd6: sine = 16'h9237;
			8'hd7: sine = 16'h93dd;
			8'hd8: sine = 16'h9594;
			8'hd9: sine = 16'h975b;
			8'hda: sine = 16'h9932;
			8'hdb: sine = 16'h9b19;
			8'hdc: sine = 16'h9d0f;
			8'hdd: sine = 16'h9f15;
			8'hde: sine = 16'ha12a;
			8'hdf: sine = 16'ha34d;
			8'he0: sine = 16'ha57f;
			8'he1: sine = 16'ha7be;
			8'he2: sine = 16'haa0c;
			8'he3: sine = 16'hac66;
			8'he4: sine = 16'haecd;
			8'he5: sine = 16'hb141;
			8'he6: sine = 16'hb3c1;
			8'he7: sine = 16'hb64d;
			8'he8: sine = 16'hb8e4;
			8'he9: sine = 16'hbb86;
			8'hea: sine = 16'hbe33;
			8'heb: sine = 16'hc0ea;
			8'hec: sine = 16'hc3aa;
			8'hed: sine = 16'hc674;
			8'hee: sine = 16'hc947;
			8'hef: sine = 16'hcc22;
			8'hf0: sine = 16'hcf05;
			8'hf1: sine = 16'hd1f0;
			8'hf2: sine = 16'hd4e2;
			8'hf3: sine = 16'hd7da;
			8'hf4: sine = 16'hdad9;
			8'hf5: sine = 16'hdddd;
			8'hf6: sine = 16'he0e7;
			8'hf7: sine = 16'he3f5;
			8'hf8: sine = 16'he708;
			8'hf9: sine = 16'hea1f;
			8'hfa: sine = 16'hed39;
			8'hfb: sine = 16'hf055;
			8'hfc: sine = 16'hf375;
			8'hfd: sine = 16'hf696;
			8'hfe: sine = 16'hf9b9;
			8'hff: sine = 16'hfcdc;
	endcase
end
endmodule

//////////////////////////////////////////////////
////////////	Square Wave ROM Table	//////////////
//////////////////////////////////////////////////
// produces a 2's comp, 16-bit, approximation
// of a square wave, given an input phase (address)
module square_rom (clock, address, square);
input clock;
input [7:0] address;
output [15:0] square;
reg signed [15:0] square;
always@(posedge clock)
begin
    case(address)
    		8'h00: square = 16'h8000;
			8'h01: square = 16'h8000;
			8'h02: square = 16'h8000;
			8'h03: square = 16'h8000;
			8'h04: square = 16'h8000;
			8'h05: square = 16'h8000;
			8'h06: square = 16'h8000;
			8'h07: square = 16'h8000;
			8'h08: square = 16'h8000;
			8'h09: square = 16'h8000;
			8'h0a: square = 16'h8000;
			8'h0b: square = 16'h8000;
			8'h0c: square = 16'h8000;
			8'h0d: square = 16'h8000;
			8'h0e: square = 16'h8000;
			8'h0f: square = 16'h8000;
			8'h10: square = 16'h8000;
			8'h11: square = 16'h8000;
			8'h12: square = 16'h8000;
			8'h13: square = 16'h8000;
			8'h14: square = 16'h8000;
			8'h15: square = 16'h8000;
			8'h16: square = 16'h8000;
			8'h17: square = 16'h8000;
			8'h18: square = 16'h8000;
			8'h19: square = 16'h8000;
			8'h1a: square = 16'h8000;
			8'h1b: square = 16'h8000;
			8'h1c: square = 16'h8000;
			8'h1d: square = 16'h8000;
			8'h1e: square = 16'h8000;
			8'h1f: square = 16'h8000;
			8'h20: square = 16'h8000;
			8'h21: square = 16'h8000;
			8'h22: square = 16'h8000;
			8'h23: square = 16'h8000;
			8'h24: square = 16'h8000;
			8'h25: square = 16'h8000;
			8'h26: square = 16'h8000;
			8'h27: square = 16'h8000;
			8'h28: square = 16'h8000;
			8'h29: square = 16'h8000;
			8'h2a: square = 16'h8000;
			8'h2b: square = 16'h8000;
			8'h2c: square = 16'h8000;
			8'h2d: square = 16'h8000;
			8'h2e: square = 16'h8000;
			8'h2f: square = 16'h8000;
			8'h30: square = 16'h8000;
			8'h31: square = 16'h8000;
			8'h32: square = 16'h8000;
			8'h33: square = 16'h8000;
			8'h34: square = 16'h8000;
			8'h35: square = 16'h8000;
			8'h36: square = 16'h8000;
			8'h37: square = 16'h8000;
			8'h38: square = 16'h8000;
			8'h39: square = 16'h8000;
			8'h3a: square = 16'h8000;
			8'h3b: square = 16'h8000;
			8'h3c: square = 16'h8000;
			8'h3d: square = 16'h8000;
			8'h3e: square = 16'h8000;
			8'h3f: square = 16'h8000;
			8'h40: square = 16'h8000;
			8'h41: square = 16'h8000;
			8'h42: square = 16'h8000;
			8'h43: square = 16'h8000;
			8'h44: square = 16'h8000;
			8'h45: square = 16'h8000;
			8'h46: square = 16'h8000;
			8'h47: square = 16'h8000;
			8'h48: square = 16'h8000;
			8'h49: square = 16'h8000;
			8'h4a: square = 16'h8000;
			8'h4b: square = 16'h8000;
			8'h4c: square = 16'h8000;
			8'h4d: square = 16'h8000;
			8'h4e: square = 16'h8000;
			8'h4f: square = 16'h8000;
			8'h50: square = 16'h8000;
			8'h51: square = 16'h8000;
			8'h52: square = 16'h8000;
			8'h53: square = 16'h8000;
			8'h54: square = 16'h8000;
			8'h55: square = 16'h8000;
			8'h56: square = 16'h8000;
			8'h57: square = 16'h8000;
			8'h58: square = 16'h8000;
			8'h59: square = 16'h8000;
			8'h5a: square = 16'h8000;
			8'h5b: square = 16'h8000;
			8'h5c: square = 16'h8000;
			8'h5d: square = 16'h8000;
			8'h5e: square = 16'h8000;
			8'h5f: square = 16'h8000;
			8'h60: square = 16'h8000;
			8'h61: square = 16'h8000;
			8'h62: square = 16'h8000;
			8'h63: square = 16'h8000;
			8'h64: square = 16'h8000;
			8'h65: square = 16'h8000;
			8'h66: square = 16'h8000;
			8'h67: square = 16'h8000;
			8'h68: square = 16'h8000;
			8'h69: square = 16'h8000;
			8'h6a: square = 16'h8000;
			8'h6b: square = 16'h8000;
			8'h6c: square = 16'h8000;
			8'h6d: square = 16'h8000;
			8'h6e: square = 16'h8000;
			8'h6f: square = 16'h8000;
			8'h70: square = 16'h8000;
			8'h71: square = 16'h8000;
			8'h72: square = 16'h8000;
			8'h73: square = 16'h8000;
			8'h74: square = 16'h8000;
			8'h75: square = 16'h8000;
			8'h76: square = 16'h8000;
			8'h77: square = 16'h8000;
			8'h78: square = 16'h8000;
			8'h79: square = 16'h8000;
			8'h7a: square = 16'h8000;
			8'h7b: square = 16'h8000;
			8'h7c: square = 16'h8000;
			8'h7d: square = 16'h8000;
			8'h7e: square = 16'h8000;
			8'h7f: square = 16'h8000;
			8'h80: square = 16'h7fff;
			8'h81: square = 16'h7fff;
			8'h82: square = 16'h7fff;
			8'h83: square = 16'h7fff;
			8'h84: square = 16'h7fff;
			8'h85: square = 16'h7fff;
			8'h86: square = 16'h7fff;
			8'h87: square = 16'h7fff;
			8'h88: square = 16'h7fff;
			8'h89: square = 16'h7fff;
			8'h8a: square = 16'h7fff;
			8'h8b: square = 16'h7fff;
			8'h8c: square = 16'h7fff;
			8'h8d: square = 16'h7fff;
			8'h8e: square = 16'h7fff;
			8'h8f: square = 16'h7fff;
			8'h90: square = 16'h7fff;
			8'h91: square = 16'h7fff;
			8'h92: square = 16'h7fff;
			8'h93: square = 16'h7fff;
			8'h94: square = 16'h7fff;
			8'h95: square = 16'h7fff;
			8'h96: square = 16'h7fff;
			8'h97: square = 16'h7fff;
			8'h98: square = 16'h7fff;
			8'h99: square = 16'h7fff;
			8'h9a: square = 16'h7fff;
			8'h9b: square = 16'h7fff;
			8'h9c: square = 16'h7fff;
			8'h9d: square = 16'h7fff;
			8'h9e: square = 16'h7fff;
			8'h9f: square = 16'h7fff;
			8'ha0: square = 16'h7fff;
			8'ha1: square = 16'h7fff;
			8'ha2: square = 16'h7fff;
			8'ha3: square = 16'h7fff;
			8'ha4: square = 16'h7fff;
			8'ha5: square = 16'h7fff;
			8'ha6: square = 16'h7fff;
			8'ha7: square = 16'h7fff;
			8'ha8: square = 16'h7fff;
			8'ha9: square = 16'h7fff;
			8'haa: square = 16'h7fff;
			8'hab: square = 16'h7fff;
			8'hac: square = 16'h7fff;
			8'had: square = 16'h7fff;
			8'hae: square = 16'h7fff;
			8'haf: square = 16'h7fff;
			8'hb0: square = 16'h7fff;
			8'hb1: square = 16'h7fff;
			8'hb2: square = 16'h7fff;
			8'hb3: square = 16'h7fff;
			8'hb4: square = 16'h7fff;
			8'hb5: square = 16'h7fff;
			8'hb6: square = 16'h7fff;
			8'hb7: square = 16'h7fff;
			8'hb8: square = 16'h7fff;
			8'hb9: square = 16'h7fff;
			8'hba: square = 16'h7fff;
			8'hbb: square = 16'h7fff;
			8'hbc: square = 16'h7fff;
			8'hbd: square = 16'h7fff;
			8'hbe: square = 16'h7fff;
			8'hbf: square = 16'h7fff;
			8'hc0: square = 16'h7fff;
			8'hc1: square = 16'h7fff;
			8'hc2: square = 16'h7fff;
			8'hc3: square = 16'h7fff;
			8'hc4: square = 16'h7fff;
			8'hc5: square = 16'h7fff;
			8'hc6: square = 16'h7fff;
			8'hc7: square = 16'h7fff;
			8'hc8: square = 16'h7fff;
			8'hc9: square = 16'h7fff;
			8'hca: square = 16'h7fff;
			8'hcb: square = 16'h7fff;
			8'hcc: square = 16'h7fff;
			8'hcd: square = 16'h7fff;
			8'hce: square = 16'h7fff;
			8'hcf: square = 16'h7fff;
			8'hd0: square = 16'h7fff;
			8'hd1: square = 16'h7fff;
			8'hd2: square = 16'h7fff;
			8'hd3: square = 16'h7fff;
			8'hd4: square = 16'h7fff;
			8'hd5: square = 16'h7fff;
			8'hd6: square = 16'h7fff;
			8'hd7: square = 16'h7fff;
			8'hd8: square = 16'h7fff;
			8'hd9: square = 16'h7fff;
			8'hda: square = 16'h7fff;
			8'hdb: square = 16'h7fff;
			8'hdc: square = 16'h7fff;
			8'hdd: square = 16'h7fff;
			8'hde: square = 16'h7fff;
			8'hdf: square = 16'h7fff;
			8'he0: square = 16'h7fff;
			8'he1: square = 16'h7fff;
			8'he2: square = 16'h7fff;
			8'he3: square = 16'h7fff;
			8'he4: square = 16'h7fff;
			8'he5: square = 16'h7fff;
			8'he6: square = 16'h7fff;
			8'he7: square = 16'h7fff;
			8'he8: square = 16'h7fff;
			8'he9: square = 16'h7fff;
			8'hea: square = 16'h7fff;
			8'heb: square = 16'h7fff;
			8'hec: square = 16'h7fff;
			8'hed: square = 16'h7fff;
			8'hee: square = 16'h7fff;
			8'hef: square = 16'h7fff;
			8'hf0: square = 16'h7fff;
			8'hf1: square = 16'h7fff;
			8'hf2: square = 16'h7fff;
			8'hf3: square = 16'h7fff;
			8'hf4: square = 16'h7fff;
			8'hf5: square = 16'h7fff;
			8'hf6: square = 16'h7fff;
			8'hf7: square = 16'h7fff;
			8'hf8: square = 16'h7fff;
			8'hf9: square = 16'h7fff;
			8'hfa: square = 16'h7fff;
			8'hfb: square = 16'h7fff;
			8'hfc: square = 16'h7fff;
			8'hfd: square = 16'h7fff;
			8'hfe: square = 16'h7fff;
			8'hff: square = 16'h7fff;
	endcase
end
endmodule

//////////////////////////////////////////////////
////////////	Saw Wave ROM Table	//////////////
//////////////////////////////////////////////////
// produces a 2's comp, 16-bit, approximation
// of a saw wave, given an input phase (address)
module saw_rom (clock, address, saw);
input clock;
input [7:0] address;
output [15:0] saw;
reg signed [15:0] saw;
always@(posedge clock)
begin
    case(address)
			8'h00: saw = 16'h7fff;
			8'h01: saw = 16'h7efe;
			8'h02: saw = 16'h7dfd;
			8'h03: saw = 16'h7cfc;
			8'h04: saw = 16'h7bfb;
			8'h05: saw = 16'h7afa;
			8'h06: saw = 16'h79f9;
			8'h07: saw = 16'h78f8;
			8'h08: saw = 16'h77f7;
			8'h09: saw = 16'h76f6;
			8'h0a: saw = 16'h75f5;
			8'h0b: saw = 16'h74f4;
			8'h0c: saw = 16'h73f3;
			8'h0d: saw = 16'h72f2;
			8'h0e: saw = 16'h71f1;
			8'h0f: saw = 16'h70f0;
			8'h10: saw = 16'h6fef;
			8'h11: saw = 16'h6eee;
			8'h12: saw = 16'h6ded;
			8'h13: saw = 16'h6cec;
			8'h14: saw = 16'h6beb;
			8'h15: saw = 16'h6aea;
			8'h16: saw = 16'h69e9;
			8'h17: saw = 16'h68e8;
			8'h18: saw = 16'h67e7;
			8'h19: saw = 16'h66e6;
			8'h1a: saw = 16'h65e5;
			8'h1b: saw = 16'h64e4;
			8'h1c: saw = 16'h63e3;
			8'h1d: saw = 16'h62e2;
			8'h1e: saw = 16'h61e1;
			8'h1f: saw = 16'h60e0;
			8'h20: saw = 16'h5fdf;
			8'h21: saw = 16'h5ede;
			8'h22: saw = 16'h5ddd;
			8'h23: saw = 16'h5cdc;
			8'h24: saw = 16'h5bdb;
			8'h25: saw = 16'h5ada;
			8'h26: saw = 16'h59d9;
			8'h27: saw = 16'h58d8;
			8'h28: saw = 16'h57d7;
			8'h29: saw = 16'h56d6;
			8'h2a: saw = 16'h55d5;
			8'h2b: saw = 16'h54d4;
			8'h2c: saw = 16'h53d3;
			8'h2d: saw = 16'h52d2;
			8'h2e: saw = 16'h51d1;
			8'h2f: saw = 16'h50d0;
			8'h30: saw = 16'h4fcf;
			8'h31: saw = 16'h4ece;
			8'h32: saw = 16'h4dcd;
			8'h33: saw = 16'h4ccc;
			8'h34: saw = 16'h4bcb;
			8'h35: saw = 16'h4aca;
			8'h36: saw = 16'h49c9;
			8'h37: saw = 16'h48c8;
			8'h38: saw = 16'h47c7;
			8'h39: saw = 16'h46c6;
			8'h3a: saw = 16'h45c5;
			8'h3b: saw = 16'h44c4;
			8'h3c: saw = 16'h43c3;
			8'h3d: saw = 16'h42c2;
			8'h3e: saw = 16'h41c1;
			8'h3f: saw = 16'h40c0;
			8'h40: saw = 16'h3fbf;
			8'h41: saw = 16'h3ebe;
			8'h42: saw = 16'h3dbd;
			8'h43: saw = 16'h3cbc;
			8'h44: saw = 16'h3bbb;
			8'h45: saw = 16'h3aba;
			8'h46: saw = 16'h39b9;
			8'h47: saw = 16'h38b8;
			8'h48: saw = 16'h37b7;
			8'h49: saw = 16'h36b6;
			8'h4a: saw = 16'h35b5;
			8'h4b: saw = 16'h34b4;
			8'h4c: saw = 16'h33b3;
			8'h4d: saw = 16'h32b2;
			8'h4e: saw = 16'h31b1;
			8'h4f: saw = 16'h30b0;
			8'h50: saw = 16'h2faf;
			8'h51: saw = 16'h2eae;
			8'h52: saw = 16'h2dad;
			8'h53: saw = 16'h2cac;
			8'h54: saw = 16'h2bab;
			8'h55: saw = 16'h2aaa;
			8'h56: saw = 16'h29a9;
			8'h57: saw = 16'h28a8;
			8'h58: saw = 16'h27a7;
			8'h59: saw = 16'h26a6;
			8'h5a: saw = 16'h25a5;
			8'h5b: saw = 16'h24a4;
			8'h5c: saw = 16'h23a3;
			8'h5d: saw = 16'h22a2;
			8'h5e: saw = 16'h21a1;
			8'h5f: saw = 16'h20a0;
			8'h60: saw = 16'h1f9f;
			8'h61: saw = 16'h1e9e;
			8'h62: saw = 16'h1d9d;
			8'h63: saw = 16'h1c9c;
			8'h64: saw = 16'h1b9b;
			8'h65: saw = 16'h1a9a;
			8'h66: saw = 16'h1999;
			8'h67: saw = 16'h1898;
			8'h68: saw = 16'h1797;
			8'h69: saw = 16'h1696;
			8'h6a: saw = 16'h1595;
			8'h6b: saw = 16'h1494;
			8'h6c: saw = 16'h1393;
			8'h6d: saw = 16'h1292;
			8'h6e: saw = 16'h1191;
			8'h6f: saw = 16'h1090;
			8'h70: saw = 16'h0f8f;
			8'h71: saw = 16'h0e8e;
			8'h72: saw = 16'h0d8d;
			8'h73: saw = 16'h0c8c;
			8'h74: saw = 16'h0b8b;
			8'h75: saw = 16'h0a8a;
			8'h76: saw = 16'h0989;
			8'h77: saw = 16'h0888;
			8'h78: saw = 16'h0787;
			8'h79: saw = 16'h0686;
			8'h7a: saw = 16'h0585;
			8'h7b: saw = 16'h0484;
			8'h7c: saw = 16'h0383;
			8'h7d: saw = 16'h0282;
			8'h7e: saw = 16'h0181;
			8'h7f: saw = 16'h0080;
			8'h80: saw = 16'hff7f;
			8'h81: saw = 16'hfe7e;
			8'h82: saw = 16'hfd7d;
			8'h83: saw = 16'hfc7c;
			8'h84: saw = 16'hfb7b;
			8'h85: saw = 16'hfa7a;
			8'h86: saw = 16'hf979;
			8'h87: saw = 16'hf878;
			8'h88: saw = 16'hf777;
			8'h89: saw = 16'hf676;
			8'h8a: saw = 16'hf575;
			8'h8b: saw = 16'hf474;
			8'h8c: saw = 16'hf373;
			8'h8d: saw = 16'hf272;
			8'h8e: saw = 16'hf171;
			8'h8f: saw = 16'hf070;
			8'h90: saw = 16'hef6f;
			8'h91: saw = 16'hee6e;
			8'h92: saw = 16'hed6d;
			8'h93: saw = 16'hec6c;
			8'h94: saw = 16'heb6b;
			8'h95: saw = 16'hea6a;
			8'h96: saw = 16'he969;
			8'h97: saw = 16'he868;
			8'h98: saw = 16'he767;
			8'h99: saw = 16'he666;
			8'h9a: saw = 16'he565;
			8'h9b: saw = 16'he464;
			8'h9c: saw = 16'he363;
			8'h9d: saw = 16'he262;
			8'h9e: saw = 16'he161;
			8'h9f: saw = 16'he060;
			8'ha0: saw = 16'hdf5f;
			8'ha1: saw = 16'hde5e;
			8'ha2: saw = 16'hdd5d;
			8'ha3: saw = 16'hdc5c;
			8'ha4: saw = 16'hdb5b;
			8'ha5: saw = 16'hda5a;
			8'ha6: saw = 16'hd959;
			8'ha7: saw = 16'hd858;
			8'ha8: saw = 16'hd757;
			8'ha9: saw = 16'hd656;
			8'haa: saw = 16'hd555;
			8'hab: saw = 16'hd454;
			8'hac: saw = 16'hd353;
			8'had: saw = 16'hd252;
			8'hae: saw = 16'hd151;
			8'haf: saw = 16'hd050;
			8'hb0: saw = 16'hcf4f;
			8'hb1: saw = 16'hce4e;
			8'hb2: saw = 16'hcd4d;
			8'hb3: saw = 16'hcc4c;
			8'hb4: saw = 16'hcb4b;
			8'hb5: saw = 16'hca4a;
			8'hb6: saw = 16'hc949;
			8'hb7: saw = 16'hc848;
			8'hb8: saw = 16'hc747;
			8'hb9: saw = 16'hc646;
			8'hba: saw = 16'hc545;
			8'hbb: saw = 16'hc444;
			8'hbc: saw = 16'hc343;
			8'hbd: saw = 16'hc242;
			8'hbe: saw = 16'hc141;
			8'hbf: saw = 16'hc040;
			8'hc0: saw = 16'hbf3f;
			8'hc1: saw = 16'hbe3e;
			8'hc2: saw = 16'hbd3d;
			8'hc3: saw = 16'hbc3c;
			8'hc4: saw = 16'hbb3b;
			8'hc5: saw = 16'hba3a;
			8'hc6: saw = 16'hb939;
			8'hc7: saw = 16'hb838;
			8'hc8: saw = 16'hb737;
			8'hc9: saw = 16'hb636;
			8'hca: saw = 16'hb535;
			8'hcb: saw = 16'hb434;
			8'hcc: saw = 16'hb333;
			8'hcd: saw = 16'hb232;
			8'hce: saw = 16'hb131;
			8'hcf: saw = 16'hb030;
			8'hd0: saw = 16'haf2f;
			8'hd1: saw = 16'hae2e;
			8'hd2: saw = 16'had2d;
			8'hd3: saw = 16'hac2c;
			8'hd4: saw = 16'hab2b;
			8'hd5: saw = 16'haa2a;
			8'hd6: saw = 16'ha929;
			8'hd7: saw = 16'ha828;
			8'hd8: saw = 16'ha727;
			8'hd9: saw = 16'ha626;
			8'hda: saw = 16'ha525;
			8'hdb: saw = 16'ha424;
			8'hdc: saw = 16'ha323;
			8'hdd: saw = 16'ha222;
			8'hde: saw = 16'ha121;
			8'hdf: saw = 16'ha020;
			8'he0: saw = 16'h9f1f;
			8'he1: saw = 16'h9e1e;
			8'he2: saw = 16'h9d1d;
			8'he3: saw = 16'h9c1c;
			8'he4: saw = 16'h9b1b;
			8'he5: saw = 16'h9a1a;
			8'he6: saw = 16'h9919;
			8'he7: saw = 16'h9818;
			8'he8: saw = 16'h9717;
			8'he9: saw = 16'h9616;
			8'hea: saw = 16'h9515;
			8'heb: saw = 16'h9414;
			8'hec: saw = 16'h9313;
			8'hed: saw = 16'h9212;
			8'hee: saw = 16'h9111;
			8'hef: saw = 16'h9010;
			8'hf0: saw = 16'h8f0f;
			8'hf1: saw = 16'h8e0e;
			8'hf2: saw = 16'h8d0d;
			8'hf3: saw = 16'h8c0c;
			8'hf4: saw = 16'h8b0b;
			8'hf5: saw = 16'h8a0a;
			8'hf6: saw = 16'h8909;
			8'hf7: saw = 16'h8808;
			8'hf8: saw = 16'h8707;
			8'hf9: saw = 16'h8606;
			8'hfa: saw = 16'h8505;
			8'hfb: saw = 16'h8404;
			8'hfc: saw = 16'h8303;
			8'hfd: saw = 16'h8202;
			8'hfe: saw = 16'h8101;
			8'hff: saw = 16'h8000;
			endcase
end
endmodule
//////////////////////////////////////////////////
